//
// CV32E40P-specific macro defintions
//
`define RISCV_CSR_MVENDORID  32'h0000_0000
`define RISCV_CSR_MARCHID  32'h0000_0000
`define RISCV_CSR_MIMPID  32'h0000_0000
`define RISCV_CSR_MHARTID  32'h0000_0000
`define RISCV_CSR_MSTATUS  32'h0000_030c
`define RISCV_CSR_MISA  32'h0000_0000
`define RISCV_CSR_MEDELEG  32'h0000_0000
`define RISCV_CSR_MIDELEG  32'h0000_0000
`define RISCV_CSR_MIE  32'h0000_0000
`define RISCV_CSR_MTVEC  32'h0000_0308
`define RISCV_CSR_MCOUNTEREN  32'h0000_0000
`define RISCV_CSR_MHPMEVENT3  32'h0000_0000
`define RISCV_CSR_MHPMEVENT4  32'h0000_0000
`define RISCV_CSR_MHPMEVENT5  32'h0000_0000
`define RISCV_CSR_MHPMEVENT6  32'h0000_0000
`define RISCV_CSR_MHPMEVENT7  32'h0000_0000
`define RISCV_CSR_MHPMEVENT8  32'h0000_0000
`define RISCV_CSR_MHPMEVENT9  32'h0000_0000
`define RISCV_CSR_MHPMEVENT10  32'h0000_0000
`define RISCV_CSR_MHPMEVENT31  32'h0000_0000
`define RISCV_CSR_MSCRATCH  32'h0000_0300
`define RISCV_CSR_MEPC  32'h0000_0310
`define RISCV_CSR_MCAUSE  32'h0000_0000
`define RISCV_CSR_MTVAL  32'h0000_0000
`define RISCV_CSR_MIP  32'h0000_0000
`define RISCV_CSR_PMPCFG0  32'h0000_0000
`define RISCV_CSR_PMPCFG2  32'h0000_0000
`define RISCV_CSR_PMPADDR0   32'h0000_0000
`define RISCV_CSR_PMPADDR1    32'h0000_0000
`define RISCV_CSR_PMPADDR2    32'h0000_0000
`define RISCV_CSR_PMPADDR3    32'h0000_0000
`define RISCV_CSR_PMPADDR4    32'h0000_0000
`define RISCV_CSR_PMPADDR5    32'h0000_0000
`define RISCV_CSR_PMPADDR6    32'h0000_0000
`define RISCV_CSR_PMPADDR7    32'h0000_0000
`define RISCV_CSR_PMPADDR8    32'h0000_0000
`define RISCV_CSR_PMPADDR9    32'h0000_0000
`define RISCV_CSR_PMPADDR10    32'h0000_0000
`define RISCV_CSR_PMPADDR11    32'h0000_0000
`define RISCV_CSR_PMPADDR12    32'h0000_0000
`define RISCV_CSR_PMPADDR13    32'h0000_0000
`define RISCV_CSR_PMPADDR14    32'h0000_0000
`define RISCV_CSR_PMPADDR15    32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER_MCYCLE  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER_MINSTRET  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER0   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER1   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER2   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER3   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER4   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER5   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER6   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER7   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER8   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER9   32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER10  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER11  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER12  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER13  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER14  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER15  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER16  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER17  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER18  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER19  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER20  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER21  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER22  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER23  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER24  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER25  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER26  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER27  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER28  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER29  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER30  32'h0000_0000
`define RISCV_CSR_MHPMCOUNTER31  32'h0000_0000
`define RISCV_CSR_MTIMECMP  32'h0000_0000
`define RISCV_CSR_SSTATUS  32'h0000_0000
`define RISCV_CSR_SIE  32'h0000_0000
`define RISCV_CSR_STVEC  32'h0000_0314
`define RISCV_CSR_SCOUNTEREN  32'h0000_0000
`define RISCV_CSR_SSCRATCH  32'h0000_0000
`define RISCV_CSR_SEPC  32'h0000_0000
`define RISCV_CSR_SCAUSE  32'h0000_0000
`define RISCV_CSR_STVAL  32'h0000_0000
`define RISCV_CSR_SIP  32'h0000_0000
`define RISCV_CSR_SATP  32'h0000_0000
`define RISCV_CSR_FFLAGS  32'h0000_0000
`define RISCV_CSR_FRM  32'h0000_0000
`define RISCV_CSR_FCSR  32'h0000_0000
`define RISCV_CSR_HPMCOUNTER_CYCLE    32'h0000_0000
`define RISCV_CSR_HPMCOUNTER_TIME     32'h0000_0000
`define RISCV_CSR_HPMCOUNTER_INSTRET  32'h0000_0000
`define RISCV_CSR_HPMCOUNTER3         32'h0000_0000
`define RISCV_CSR_HPMCOUNTER4         32'h0000_0000
`define RISCV_CSR_HPMCOUNTER5         32'h0000_0000
`define RISCV_CSR_HPMCOUNTER6         32'h0000_0000
`define RISCV_CSR_HPMCOUNTER7         32'h0000_0000
`define RISCV_CSR_HPMCOUNTER8         32'h0000_0000
`define RISCV_CSR_HPMCOUNTER9         32'h0000_0000
`define RISCV_CSR_HPMCOUNTER10        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER11        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER12        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER13        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER14        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER15        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER16        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER17        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER18        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER19        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER20        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER21        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER22        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER23        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER24        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER25        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER26        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER27        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER28        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER29        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER30        32'h0000_0000
`define RISCV_CSR_HPMCOUNTER31        32'h0000_0000

`define RISCV_CSR_PMPCFG0_PMP7A_OFF   32'h0000_0000
`define RISCV_CSR_PMPCFG0_PMP7A_TOR   32'h0000_0000
`define RISCV_CSR_PMPCFG0_PMP7A_NA4   32'h0000_0000
`define RISCV_CSR_PMPCFG0_PMP7A_NAPOT 32'h0000_0000

// These should be defined elsewhere, but are not.
// Setting to 'h0 just for compile-time tests.
`define CSR_TSELECT      32'h0000_0000
`define CSR_TDATA1       32'h0000_0000
`define CSR_TDATA2       32'h0000_0000
`define CSR_DCSR         32'h0000_0000
`define CSR_TSELECT      32'h0000_0000
`define CSR_TDATA1       32'h0000_0000
`define CSR_TDATA2       32'h0000_0000
`define CSR_DCSR         32'h0000_0000
`define CSR_TSELECT      32'h0000_0000
`define CSR_TDATA1       32'h0000_0000
`define CSR_TDATA2       32'h0000_0000
`define CSR_DCSR         32'h0000_0000
`define CSR_MSCRATCH2    32'h0000_0304
`define CSR_SSCRATCH2    32'h0000_0000
 
